* uA741 operational amplifier

.width out=80 

vcc 27 0  15.0
vee 26 0 -15.0
*vin 30 0 dc 0
vin 30 0 pulse 0 1 1e-8 1e-9
*cl 24 0 1p

rs1 1 30 1k
*rs2 2 31 1k
rs2 2 24 1k
rf 24 1 100k
r1 10 26 1k
r2 9 26 50k
r3 11 26 1k
r4 12 26 3k
r5 15 17 39k
r6 21 20 40k
r7 14 26 50k
r8 18 26 50.0
r9 24 25 25.0
r10 23 24 50.0
r11 13 26 50k
cc 22 8 30p
q1 3 2 4 qnl
q2 3 1 5 qnl
q3 7 6 4 qpl
q4 8 6 5 qpl
q5 7 9 10 qnl
q6 8 9 11 qnl
q7 27 7 9 qnl
q8 6 15 12 qnl
q9 15 15 26 qnl
q10 3 3 27 qpl
q11 6 3 27 qpl
q12 17 17 27 qpl
q13 8 13 26 qnl
q14 22 17 27 qpl
q15 22 22 21 qnl
q16 22 21 20 qnl
q17 13 13 26 qnl
q18 27 8 14 qnl
q19 20 14 18 qnl
q20 22 23 24 qnl
q21 13 25 24 qpl
q22 27 22 23 qnl
q23 26 20 25 qpl
.model qnl npn(bf=80 rb=0 cje=3p cjc=2p va=50)
.model qpl pnp(bf=10 rb=0 cje=6p cjc=4p va=50)

.op

*.plot dc v(2)
*.dc vin -1 1 0.01

*.plot ac vdb(2) vp(2)
*.ac dec 20 1 10meg

.plot tran v(1) v(2)
*.plot tran v(2)
*.tran 2.5u 250u
.tran 1e-9 1e-7

.end
